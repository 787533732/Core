`include "../core/define.v"
module exec 
(
    input   wire                    clk_i                   ,
    input   wire                    rstn_i                   ,
    //hazard detect无延迟给到E1的数据
    input   wire                    opcode_valid_i          ,
    input   wire [31:0]             opcode_opcode_i         ,
    input   wire [31:0]             opcode_pc_i             ,
    input   wire                    opcode_invalid_i        ,
    input   wire [ 4:0]             opcode_rd_idx_i         ,
    input   wire [ 4:0]             opcode_ra_idx_i         ,
    input   wire [ 4:0]             opcode_rb_idx_i         ,
    input   wire [31:0]             opcode_ra_operand_i     ,
    input   wire [31:0]             opcode_rb_operand_i     , 
    input   wire                    hold_i                  ,
    //都是组合逻辑打一拍输出
    output  wire [31:0]             writeback_value_o       ,
    output  wire                    branch_request_o        ,//分支指令标志
    output  wire                    branch_is_taken_o       ,    
    output  wire                    branch_is_not_taken_o   ,
    output  wire [31:0]             branch_pc_o             ,          
    output  wire [31:0]             branch_source_o         ,      
    output  wire                    branch_call_o           ,        
    output  wire                    branch_ret_o            ,         
    output  wire                    branch_jmp_o            ,
    //组合逻辑的输出，没有打一拍    
    output  wire                    branch_d_request_o      ,
    output  wire [31:0]             branch_d_pc_o           ,
    output  wire [ 1:0]             branch_d_priv_o          
);   
//-------------------------------------------------------------
//立即数拓展
//-------------------------------------------------------------
    wire [31:0] imm20_w  = {opcode_opcode_i[31:12], 12'b0};//LUI，AUIPC
    wire [31:0] imm12_w  = {{20{opcode_opcode_i[31]}}, opcode_opcode_i[31:20]};
    wire [31:0] bimm_w   = {{20{opcode_opcode_i[31]}}, opcode_opcode_i[7], opcode_opcode_i[30:25], opcode_opcode_i[11:8], 1'b0};//B-Type
    wire [31:0] jimm20_w = {{12{opcode_opcode_i[31]}}, opcode_opcode_i[19:12], opcode_opcode_i[20], opcode_opcode_i[30:21], 1'b0};//JAL
    wire [ 4:0] shamt_w  = opcode_opcode_i[24:20];

//-------------------------------------------------------------
//算术逻辑操作
//-------------------------------------------------------------
    reg [ 3:0] alu_func_r;
    reg [31:0] alu_input_a_r;
    reg [31:0] alu_input_b_r;

    always @(*) begin
        alu_func_r    = `ALU_NONE;
        alu_input_a_r = 32'h0;
        alu_input_b_r = 32'h0;       
        if     ((opcode_opcode_i & `INST_ADD_MASK) == `INST_ADD) begin//1ADD
            alu_func_r    = `ALU_ADD;
            alu_input_a_r = opcode_ra_operand_i;
            alu_input_b_r = opcode_rb_operand_i;     
        end
        else if((opcode_opcode_i & `INST_SUB_MASK) == `INST_SUB) begin//2SUB
            alu_func_r     = `ALU_SUB;
            alu_input_a_r  = opcode_ra_operand_i;
            alu_input_b_r  = opcode_rb_operand_i;
        end
        else if((opcode_opcode_i & `INST_SLL_MASK) == `INST_SLL) begin//3SLL
            alu_func_r     = `ALU_SHIFTL;
            alu_input_a_r  = opcode_ra_operand_i;
            alu_input_b_r  = opcode_rb_operand_i;
        end
        else if((opcode_opcode_i & `INST_SLT_MASK) == `INST_SLT) begin//4SLT
            alu_func_r     = `ALU_LESS_THAN_SIGNED;
            alu_input_a_r  = opcode_ra_operand_i;
            alu_input_b_r  = opcode_rb_operand_i;
        end
        else if((opcode_opcode_i & `INST_SLTU_MASK) == `INST_SLTU) begin//5SLTU
            alu_func_r     = `ALU_LESS_THAN;
            alu_input_a_r  = opcode_ra_operand_i;
            alu_input_b_r  = opcode_rb_operand_i;
        end
        else if((opcode_opcode_i & `INST_XOR_MASK) == `INST_XOR) begin//6XOR
            alu_func_r     = `ALU_XOR;
            alu_input_a_r  = opcode_ra_operand_i;
            alu_input_b_r  = opcode_rb_operand_i;
        end
        else if((opcode_opcode_i & `INST_SRL_MASK) == `INST_SRL) begin//7SRL
            alu_func_r     = `ALU_SHIFTR;
            alu_input_a_r  = opcode_ra_operand_i;
            alu_input_b_r  = opcode_rb_operand_i;
        end
        else if((opcode_opcode_i & `INST_SRA_MASK) == `INST_SRA) begin//8SRA
            alu_func_r     = `ALU_SHIFTR_ARITH;
            alu_input_a_r  = opcode_ra_operand_i;
            alu_input_b_r  = opcode_rb_operand_i;
        end
        else if((opcode_opcode_i & `INST_OR_MASK) == `INST_OR) begin//9OR
            alu_func_r     = `ALU_OR;
            alu_input_a_r  = opcode_ra_operand_i;
            alu_input_b_r  = opcode_rb_operand_i;
        end
        else if((opcode_opcode_i & `INST_AND_MASK) == `INST_AND) begin//10AND
            alu_func_r     = `ALU_AND;
            alu_input_a_r  = opcode_ra_operand_i;
            alu_input_b_r  = opcode_rb_operand_i;
        end
        else if((opcode_opcode_i & `INST_ADDI_MASK) == `INST_ADDI) begin//11ADDI
            alu_func_r     = `ALU_ADD;
            alu_input_a_r  = opcode_ra_operand_i;
            alu_input_b_r  = imm12_w;
        end
        else if((opcode_opcode_i & `INST_SLTI_MASK) == `INST_SLTI) begin//12SLTI
            alu_func_r     = `ALU_LESS_THAN_SIGNED;
            alu_input_a_r  = opcode_ra_operand_i;
            alu_input_b_r  = imm12_w;
        end
        else if((opcode_opcode_i & `INST_SLTIU_MASK) == `INST_SLTIU) begin//13SLTIU
            alu_func_r     = `ALU_LESS_THAN;
            alu_input_a_r  = opcode_ra_operand_i;
            alu_input_b_r  = imm12_w;
        end
        else if((opcode_opcode_i & `INST_XORI_MASK) == `INST_XORI) begin//14XORI
            alu_func_r     = `ALU_XOR;
            alu_input_a_r  = opcode_ra_operand_i;
            alu_input_b_r  = imm12_w;
        end
        else if((opcode_opcode_i & `INST_ORI_MASK) == `INST_ORI) begin//15ORI
            alu_func_r     = `ALU_OR;
            alu_input_a_r  = opcode_ra_operand_i;
            alu_input_b_r  = imm12_w;
        end
        else if((opcode_opcode_i & `INST_ANDI_MASK) == `INST_ANDI) begin//16ANDI
            alu_func_r     = `ALU_AND;
            alu_input_a_r  = opcode_ra_operand_i;
            alu_input_b_r  = imm12_w;
        end
        else if((opcode_opcode_i & `INST_SLLI_MASK) == `INST_SLLI) begin//17SLLI
            alu_func_r     = `ALU_SHIFTL;
            alu_input_a_r  = opcode_ra_operand_i;
            alu_input_b_r  = {27'b0, shamt_w};
        end
        else if((opcode_opcode_i & `INST_SRLI_MASK) == `INST_SRLI) begin//18SRLI
            alu_func_r     = `ALU_SHIFTR;
            alu_input_a_r  = opcode_ra_operand_i;
            alu_input_b_r  = {27'b0, shamt_w};
        end
        else if((opcode_opcode_i & `INST_SRAI_MASK) == `INST_SRAI) begin//19SRAI
            alu_func_r     = `ALU_SHIFTR_ARITH;
            alu_input_a_r  = opcode_ra_operand_i;
            alu_input_b_r  = {27'b0, shamt_w};
        end
        else if((opcode_opcode_i & `INST_LUI_MASK) == `INST_LUI) begin//20LUI
            alu_input_a_r  = imm20_w;
        end
        else if((opcode_opcode_i & `INST_AUIPC_MASK) == `INST_AUIPC) begin//21AUIPC
            alu_func_r     = `ALU_ADD;
            alu_input_a_r  = opcode_pc_i;
            alu_input_b_r  = imm20_w;
        end     
        else if(((opcode_opcode_i & `INST_JAL_MASK) == `INST_JAL) || ((opcode_opcode_i & `INST_JALR_MASK) == `INST_JALR)) begin//22JAL,23JALR
            alu_func_r     = `ALU_ADD;
            alu_input_a_r  = opcode_pc_i;
            alu_input_b_r  = 32'd4;
        end
    end    

    wire [31:0] alu_p_w;
    alu u_alu
    (
        .alu_op_i           (alu_func_r   ),
        .alu_a_i            (alu_input_a_r),
        .alu_b_i            (alu_input_b_r),

        .alu_p_o            (alu_p_w      )
    );
    //ALU输出打一拍
    reg [31:0] result_q;
    always @(posedge clk_i or negedge rstn_i) begin
        if(!rstn_i)
            result_q <= 32'h0;
        else if(~hold_i)
            result_q <= alu_p_w;
    end
    assign writeback_value_o = result_q;
//-------------------------------------------------------------
// 定义两个比大小的函数
//-------------------------------------------------------------
    //如果x<y(signed)输出1
    function [0:0] less_than_signed;
    input  [31:0] x;
    input  [31:0] y;
    reg [31:0] v;
    begin
        v = (x - y); 
        if (x[31] != y[31])
            less_than_signed = x[31];
        else
            less_than_signed = v[31];
    end
    endfunction
    //如果x>y(signed)输出1
    function [0:0] greater_than_signed;
        input  [31:0] x;
        input  [31:0] y;
        reg [31:0] v;
    begin
        v = (y - x); 
        if (x[31] != y[31]) 
            greater_than_signed = y[31];
        else
            greater_than_signed = v[31];
    end
    endfunction

//-------------------------------------------------------------
// Execute 分支跳转判断
//------------------------------------------------------------
    reg         branch_r;
    reg         branch_taken_r;
    reg [31:0]  branch_target_r;
    reg         branch_call_r;
    reg         branch_ret_r; 
    reg         branch_jmp_r; 
    always @(*) begin
        branch_r        = 1'b0;
        branch_taken_r  = 1'b0;
        branch_target_r = opcode_pc_i + bimm_w;//默认B型指令的跳转地址
        //call ret jmp暂不了解
        branch_call_r   = 1'b0;
        branch_ret_r    = 1'b0;
        branch_jmp_r    = 1'b0;
        if     ((opcode_opcode_i & `INST_BEQ_MASK) == `INST_BEQ) begin//1BEQ
            branch_r       = 1'b1;
            branch_taken_r = (opcode_ra_operand_i == opcode_rb_operand_i);
        end
        else if((opcode_opcode_i & `INST_BNE_MASK) == `INST_BNE) begin//2BNE
            branch_r       = 1'b1;    
            branch_taken_r = (opcode_ra_operand_i != opcode_rb_operand_i);
        end
        else if((opcode_opcode_i & `INST_BLT_MASK) == `INST_BLT) begin//3BLT
    
            branch_r       = 1'b1;
            branch_taken_r = less_than_signed(opcode_ra_operand_i, opcode_rb_operand_i);
        end
        else if((opcode_opcode_i & `INST_BGE_MASK) == `INST_BGE) begin//4BGE
            branch_r       = 1'b1;    
            branch_taken_r = greater_than_signed(opcode_ra_operand_i,opcode_rb_operand_i) | (opcode_ra_operand_i == opcode_rb_operand_i);
        end
        else if((opcode_opcode_i & `INST_BLTU_MASK) == `INST_BLTU) begin//5BLTU
            branch_r       = 1'b1;    
            branch_taken_r = (opcode_ra_operand_i < opcode_rb_operand_i);
        end
        else if((opcode_opcode_i & `INST_BGEU_MASK) == `INST_BGEU) begin//6BGEU
            branch_r       = 1'b1;
            branch_taken_r = (opcode_ra_operand_i >= opcode_rb_operand_i);
        end 
        else if((opcode_opcode_i & `INST_JAL_MASK) == `INST_JAL) begin// jal
            branch_r        = 1'b1;
            branch_taken_r  = 1'b1;
            branch_target_r = opcode_pc_i + jimm20_w;
            branch_call_r   = (opcode_rd_idx_i == 5'd1); // RA
            branch_jmp_r    = 1'b1;
        end
        else if((opcode_opcode_i & `INST_JALR_MASK) == `INST_JALR) begin// jalr
            branch_r            = 1'b1;
            branch_taken_r      = 1'b1;
            branch_target_r     = opcode_ra_operand_i + imm12_w;
            branch_target_r[0]  = 1'b0;
            branch_ret_r        = (opcode_ra_idx_i == 5'd1 && imm12_w[11:0] == 12'b0); // RA
            branch_call_r       = !branch_ret_r && (opcode_rd_idx_i == 5'd1); // RA
            branch_jmp_r        = !branch_call_r && !branch_ret_r;
        end
    end
    //打一拍
    reg         branch_taken_q;
    reg         branch_ntaken_q;
    reg [31:0]  next_pc_q;
    reg [31:0]  current_pc_q;
    reg         branch_call_q;
    reg         branch_ret_q;
    reg         branch_jmp_q;

    always @(posedge clk_i or negedge rstn_i) begin
        if(!rstn_i) begin
            branch_taken_q  <= 1'b0;    
            branch_ntaken_q <= 1'b0;     
            next_pc_q       <= 32'h0;
            current_pc_q    <= 32'h0;  
            branch_call_q   <= 1'b0;   
            branch_ret_q    <= 1'b0;  
            branch_jmp_q    <= 1'b0; 
        end
        else if(opcode_valid_i) begin
            branch_taken_q  <= opcode_valid_i && branch_r && branch_taken_r;
            branch_ntaken_q <= opcode_valid_i && branch_r && ~branch_taken_r;
            next_pc_q       <= branch_taken_r ? branch_target_r : opcode_pc_i + 32'd4;
            current_pc_q    <= opcode_pc_i;
            branch_call_q   <= opcode_valid_i && branch_r && branch_call_r;
            branch_ret_q    <= opcode_valid_i && branch_r && branch_ret_r;
            branch_jmp_q    <= opcode_valid_i && branch_r && branch_jmp_r;
        end
    end
    //产生分支预测学习信号
    assign branch_request_o      = branch_taken_q | branch_ntaken_q;//分支指令标志
    assign branch_is_taken_o     = branch_taken_q;
    assign branch_is_not_taken_o = branch_ntaken_q;
    assign branch_pc_o           = next_pc_q;
    assign branch_source_o       = current_pc_q;
    assign branch_call_o         = branch_call_q;
    assign branch_ret_o          = branch_ret_q;
    assign branch_jmp_o          = branch_jmp_q;
    //组合逻辑的输出，没有打一拍
    assign branch_d_request_o = (branch_r && opcode_valid_i && branch_taken_r);
    assign branch_d_pc_o      = branch_target_r;
    assign branch_d_priv_o    = 2'b0; // don't care
endmodule